library IEEE;
use IEEE.std_logic_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity shifter is
port(
	I     : in std_logic;
	T     : in std_logic_vector(1 downto 0);
	Cs    : in std_logic_vector(4 downto 0);
	var   : in std_logic_vector(31 downto 0);
	Sout  : out std_logic_vector(31 downto 0)
	);
end shifter;

architecture beh of shifter is

signal v1     : std_logic_vector(31 downto 0) := X"00000000";
begin
	
	process(I,T,Cs,var)
	begin	
		if(I = '0') then
			
				if(T = "00" ) then
					if(Cs ="00000") then
						v1 <= var;
					elsif(Cs ="00001") then
						v1 <=  std_logic_vector(unsigned(var) sll 1);
					elsif(Cs = "00010") then
						v1 <=  std_logic_vector(unsigned(var) sll 2);
					elsif(Cs = "00011") then
						v1 <=  std_logic_vector(unsigned(var) sll 3);
					elsif(Cs = "00100") then
						v1 <=  std_logic_vector(unsigned(var) sll 4);
					elsif(Cs = "00101") then
						v1 <=  std_logic_vector(unsigned(var) sll 5);
					elsif(Cs = "00101") then
						v1 <=  std_logic_vector(unsigned(var) sll 6);
					elsif(Cs = "00110") then
						v1 <=  std_logic_vector(unsigned(var) sll 7);
					elsif(Cs = "00111") then
						v1 <=  std_logic_vector(unsigned(var) sll 8);
					elsif(Cs = "01000") then
						v1 <=  std_logic_vector(unsigned(var) sll 9);
					elsif(Cs = "01001") then
						v1 <=  std_logic_vector(unsigned(var) sll 10);
					elsif(Cs = "01010") then
						v1 <=  std_logic_vector(unsigned(var) sll 11);
					elsif(Cs = "01011") then
						v1 <=  std_logic_vector(unsigned(var) sll 12);
					elsif(Cs = "01100") then
						v1 <=  std_logic_vector(unsigned(var) sll 13);
					elsif(Cs = "01101") then
						v1 <=  std_logic_vector(unsigned(var) sll 14);
					elsif(Cs = "01110") then
						v1 <=  std_logic_vector(unsigned(var) sll 15);
					elsif(Cs = "01111") then
						v1 <=  std_logic_vector(unsigned(var) sll 16);
					elsif(Cs = "10000") then
						v1 <=  std_logic_vector(unsigned(var) sll 17);
					elsif(Cs = "10001") then
						v1 <=  std_logic_vector(unsigned(var) sll 18);
					elsif(Cs = "10010") then
						v1 <=  std_logic_vector(unsigned(var) sll 19);
					elsif(Cs = "10011") then
						v1 <=  std_logic_vector(unsigned(var) sll 20);
					elsif(Cs = "10100") then
						v1 <=  std_logic_vector(unsigned(var) sll 21);
					elsif(Cs = "10101") then
						v1 <=  std_logic_vector(unsigned(var) sll 22);
					elsif(Cs = "10110") then
						v1 <=  std_logic_vector(unsigned(var) sll 23);
					elsif(Cs = "10111") then
						v1 <=  std_logic_vector(unsigned(var) sll 24);
					elsif(Cs = "11000") then
						v1 <=  std_logic_vector(unsigned(var) sll 25);
					elsif(Cs = "11001") then
						v1 <=  std_logic_vector(unsigned(var) sll 25);
					elsif(Cs = "11010") then
						v1 <=  std_logic_vector(unsigned(var) sll 26);
					elsif(Cs = "11011") then
						v1 <=  std_logic_vector(unsigned(var) sll 27);
					elsif(Cs = "11100") then
						v1 <=  std_logic_vector(unsigned(var) sll 28);
					elsif(Cs = "11101") then
						v1 <=  std_logic_vector(unsigned(var) sll 29);
					elsif(Cs = "11110") then
						v1 <=  std_logic_vector(unsigned(var) sll 30);
					elsif(Cs = "11111") then
						v1 <=  std_logic_vector(unsigned(var) sll 31);
					end if;
				elsif(T = "01" ) then
					if(Cs ="00000") then
						v1 <= var;
					elsif(Cs ="00001") then
						v1 <=  std_logic_vector(unsigned(var) srl 1);
					elsif(Cs = "00010") then
						v1 <=  std_logic_vector(unsigned(var) srl 2);
					elsif(Cs = "00011") then
						v1 <=  std_logic_vector(unsigned(var) srl 3);
					elsif(Cs = "00100") then
						v1 <=  std_logic_vector(unsigned(var) srl 4);
					elsif(Cs = "00101") then
						v1 <=  std_logic_vector(unsigned(var) srl 5);
					elsif(Cs = "00101") then
						v1 <=  std_logic_vector(unsigned(var) srl 6);
					elsif(Cs = "00110") then
						v1 <=  std_logic_vector(unsigned(var) srl 7);
					elsif(Cs = "00111") then
						v1 <=  std_logic_vector(unsigned(var) srl 8);
					elsif(Cs = "01000") then
						v1 <=  std_logic_vector(unsigned(var) srl 9);
					elsif(Cs = "01001") then
						v1 <=  std_logic_vector(unsigned(var) srl 10);
					elsif(Cs = "01010") then
						v1 <=  std_logic_vector(unsigned(var) srl 11);
					elsif(Cs = "01011") then
						v1 <=  std_logic_vector(unsigned(var) srl 12);
					elsif(Cs = "01100") then
						v1 <=  std_logic_vector(unsigned(var) srl 13);
					elsif(Cs = "01101") then
						v1 <=  std_logic_vector(unsigned(var) srl 14);
					elsif(Cs = "01110") then
						v1 <=  std_logic_vector(unsigned(var) srl 15);
					elsif(Cs = "01111") then
						v1 <=  std_logic_vector(unsigned(var) srl 16);
					elsif(Cs = "10000") then
						v1 <=  std_logic_vector(unsigned(var) srl 17);
					elsif(Cs = "10001") then
						v1 <=  std_logic_vector(unsigned(var) srl 18);
					elsif(Cs = "10010") then
						v1 <=  std_logic_vector(unsigned(var) srl 19);
					elsif(Cs = "10011") then
						v1 <=  std_logic_vector(unsigned(var) srl 20);
					elsif(Cs = "10100") then
						v1 <=  std_logic_vector(unsigned(var) srl 21);
					elsif(Cs = "10101") then
						v1 <=  std_logic_vector(unsigned(var) srl 22);
					elsif(Cs = "10110") then
						v1 <=  std_logic_vector(unsigned(var) srl 23);
					elsif(Cs = "10111") then
						v1 <=  std_logic_vector(unsigned(var) srl 24);
					elsif(Cs = "11000") then
						v1 <=  std_logic_vector(unsigned(var) srl 25);
					elsif(Cs = "11001") then
						v1 <=  std_logic_vector(unsigned(var) srl 25);
					elsif(Cs = "11010") then
						v1 <=  std_logic_vector(unsigned(var) srl 26);
					elsif(Cs = "11011") then
						v1 <=  std_logic_vector(unsigned(var) srl 27);
					elsif(Cs = "11100") then
						v1 <=  std_logic_vector(unsigned(var) srl 28);
					elsif(Cs = "11101") then
						v1 <=  std_logic_vector(unsigned(var) srl 29);
					elsif(Cs = "11110") then
						v1 <=  std_logic_vector(unsigned(var) srl 30);
					elsif(Cs = "11111") then
						v1 <=  std_logic_vector(unsigned(var) srl 31);
					end if;
				elsif(T = "10" ) then
					if(Cs ="00000") then
						v1 <= var;
					elsif(Cs ="00001") then
						v1 <= var(31) & var(31 downto 1) ;
					elsif(Cs = "00010") then
						v1 <= var(31) & var(31)  & var(31 downto 2) ;
					elsif(Cs = "00011") then
						v1 <= var(31) &var(31) &var(31)  & var(31 downto 3) ;
					elsif(Cs = "00100") then
						v1 <= var(31) &var(31) &var(31)  & var(31) & var(31 downto 4) ;
					elsif(Cs = "00101") then
						v1 <= var(31) &var(31) &var(31)  & var(31) & var(31) & var(31 downto 5) ;
					elsif(Cs = "00101") then
						v1 <= var(31) &var(31) &var(31)  & var(31) & var(31) & var(31) & var(31 downto 6) ;
					elsif(Cs = "00110") then
						v1 <= var(31) &var(31) &var(31)  & var(31) & var(31) & var(31) & var(31) & var(31 downto 7) ;
					elsif(Cs = "00111") then
						v1 <=var(31) &var(31) &var(31)  & var(31) & var(31) & var(31) & var(31) & var(31) & var(31 downto 8) ;
					elsif(Cs = "01000") then
						v1 <= var(31) &var(31) &var(31)  & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31 downto 9) ;
					elsif(Cs = "01001") then
						v1 <= var(31) &var(31) &var(31)  & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31 downto 10) ;
					elsif(Cs = "01010") then
						v1 <= var(31) &var(31) &var(31)  & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31 downto 11) ;
					elsif(Cs = "01011") then
						v1 <= var(31) &var(31) &var(31)  & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31 downto 12) ;
					elsif(Cs = "01100") then
						v1 <= var(31) &var(31) &var(31)  & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31 downto 13) ;
					elsif(Cs = "01101") then
						v1 <= var(31) &var(31) &var(31)  & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31 downto 14) ;
					elsif(Cs = "01110") then
						v1 <= var(31) &var(31) &var(31)  & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31 downto 15) ;
					elsif(Cs = "01111") then
						v1 <= var(31) &var(31) &var(31)  & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31 downto 16) ;
					elsif(Cs = "10000") then
						v1 <= var(31) &var(31) &var(31)  & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31 downto 17);
					elsif(Cs = "10001") then
						v1 <= var(31) &var(31) &var(31)  & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31 downto 18) ;
					elsif(Cs = "10010") then
						v1 <= var(31) &var(31) &var(31)  & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31 downto 19) ;
					elsif(Cs = "10011") then
						v1 <= var(31) &var(31) &var(31)  & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31 downto 20) ;
					elsif(Cs = "10100") then
						v1 <= var(31) &var(31) &var(31)  & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31 downto 21) ;
					elsif(Cs = "10101") then
						v1 <= var(31) &var(31) &var(31)  & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31 downto 22) ;
					elsif(Cs = "10110") then
						v1 <= var(31) &var(31) &var(31)  & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31 downto 23) ;
					elsif(Cs = "10111") then
						v1 <= var(31) &var(31) &var(31)  & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31 downto 24) ;
					elsif(Cs = "11000") then
						v1 <= var(31) &var(31) &var(31)  & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31 downto 25) ;
					elsif(Cs = "11001") then
						v1 <= var(31) &var(31) &var(31)  & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31 downto 26) ;
					elsif(Cs = "11010") then
						v1 <= var(31) &var(31) &var(31)  & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31 downto 27);	
					elsif(Cs = "11011") then
						v1 <= var(31) &var(31) &var(31)  & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31 downto 28) ;
					elsif(Cs = "11100") then
						v1 <= var(31) &var(31) &var(31)  & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31 downto 29) ;
					elsif(Cs = "11101") then
						v1 <= var(31) &var(31) &var(31)  & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31 downto 30) ;
					elsif(Cs = "11110") then
						v1 <= var(31) &var(31) &var(31)  & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) ;
					elsif(Cs = "11111") then
						v1 <= var(31) &var(31) &var(31)  & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) & var(31) ;
					end if;
				elsif(T = "11" ) then
					if(Cs ="00000") then
						v1 <= var;
					elsif(Cs ="00001") then
						v1 <=  std_logic_vector(unsigned(var) ror 1);
					elsif(Cs = "00010") then
						v1 <=  std_logic_vector(unsigned(var) ror 2);
					elsif(Cs = "00011") then
						v1 <=  std_logic_vector(unsigned(var) ror 3);
					elsif(Cs = "00100") then
						v1 <=  std_logic_vector(unsigned(var) ror 4);
					elsif(Cs = "00101") then
						v1 <=  std_logic_vector(unsigned(var) ror 5);
					elsif(Cs = "00101") then
						v1 <=  std_logic_vector(unsigned(var) ror 6);
					elsif(Cs = "00110") then
						v1 <=  std_logic_vector(unsigned(var) ror 7);
					elsif(Cs = "00111") then
						v1 <=  std_logic_vector(unsigned(var) ror 8);
					elsif(Cs = "01000") then
						v1 <=  std_logic_vector(unsigned(var) ror 9);
					elsif(Cs = "01001") then
						v1 <=  std_logic_vector(unsigned(var) ror 10);
					elsif(Cs = "01010") then
						v1 <=  std_logic_vector(unsigned(var) ror 11);
					elsif(Cs = "01011") then
						v1 <=  std_logic_vector(unsigned(var) ror 12);
					elsif(Cs = "01100") then
						v1 <=  std_logic_vector(unsigned(var) ror 13);
					elsif(Cs = "01101") then
						v1 <=  std_logic_vector(unsigned(var) ror 14);
					elsif(Cs = "01110") then
						v1 <=  std_logic_vector(unsigned(var) ror 15);
					elsif(Cs = "01111") then
						v1 <=  std_logic_vector(unsigned(var) ror 16);
					elsif(Cs = "10000") then
						v1 <=  std_logic_vector(unsigned(var) ror 17);
					elsif(Cs = "10001") then
						v1 <=  std_logic_vector(unsigned(var) ror 18);
					elsif(Cs = "10010") then
						v1 <=  std_logic_vector(unsigned(var) ror 19);
					elsif(Cs = "10011") then
						v1 <=  std_logic_vector(unsigned(var) ror 20);
					elsif(Cs = "10100") then
						v1 <=  std_logic_vector(unsigned(var) ror 21);
					elsif(Cs = "10101") then
						v1 <=  std_logic_vector(unsigned(var) ror 22);
					elsif(Cs = "10110") then
						v1 <=  std_logic_vector(unsigned(var) ror 23);
					elsif(Cs = "10111") then
						v1 <=  std_logic_vector(unsigned(var) ror 24);
					elsif(Cs = "11000") then
						v1 <=  std_logic_vector(unsigned(var) ror 25);
					elsif(Cs = "11001") then
						v1 <=  std_logic_vector(unsigned(var) ror 25);
					elsif(Cs = "11010") then
						v1 <=  std_logic_vector(unsigned(var) ror 26);
					elsif(Cs = "11011") then
						v1 <=  std_logic_vector(unsigned(var) ror 27);
					elsif(Cs = "11100") then
						v1 <=  std_logic_vector(unsigned(var) ror 28);
					elsif(Cs = "11101") then
						v1 <=  std_logic_vector(unsigned(var) ror 29);
					elsif(Cs = "11110") then
						v1 <=  std_logic_vector(unsigned(var) ror 30);
					elsif(Cs = "11111") then
						v1 <=  std_logic_vector(unsigned(var) ror 31);
					end if;
				end if;
			elsif( I = '1') then
					if(Cs ="00000") then
						v1 <= var;
					elsif(Cs ="00001") then
						v1 <=  std_logic_vector(unsigned(var) ror 1);
					elsif(Cs = "00010") then
						v1 <=  std_logic_vector(unsigned(var) ror 2);
					elsif(Cs = "00011") then
						v1 <=  std_logic_vector(unsigned(var) ror 3);
					elsif(Cs = "00100") then
						v1 <=  std_logic_vector(unsigned(var) ror 4);
					elsif(Cs = "00101") then
						v1 <=  std_logic_vector(unsigned(var) ror 5);
					elsif(Cs = "00101") then
						v1 <=  std_logic_vector(unsigned(var) ror 6);
					elsif(Cs = "00110") then
						v1 <=  std_logic_vector(unsigned(var) ror 7);
					elsif(Cs = "00111") then
						v1 <=  std_logic_vector(unsigned(var) ror 8);
					elsif(Cs = "01000") then
						v1 <=  std_logic_vector(unsigned(var) ror 9);
					elsif(Cs = "01001") then
						v1 <=  std_logic_vector(unsigned(var) ror 10);
					elsif(Cs = "01010") then
						v1 <=  std_logic_vector(unsigned(var) ror 11);
					elsif(Cs = "01011") then
						v1 <=  std_logic_vector(unsigned(var) ror 12);
					elsif(Cs = "01100") then
						v1 <=  std_logic_vector(unsigned(var) ror 13);
					elsif(Cs = "01101") then
						v1 <=  std_logic_vector(unsigned(var) ror 14);
					elsif(Cs = "01110") then
						v1 <=  std_logic_vector(unsigned(var) ror 15);
					elsif(Cs = "01111") then
						v1 <=  std_logic_vector(unsigned(var) ror 16);
					elsif(Cs = "10000") then
						v1 <=  std_logic_vector(unsigned(var) ror 17);
					elsif(Cs = "10001") then
						v1 <=  std_logic_vector(unsigned(var) ror 18);
					elsif(Cs = "10010") then
						v1 <=  std_logic_vector(unsigned(var) ror 19);
					elsif(Cs = "10011") then
						v1 <=  std_logic_vector(unsigned(var) ror 20);
					elsif(Cs = "10100") then
						v1 <=  std_logic_vector(unsigned(var) ror 21);
					elsif(Cs = "10101") then
						v1 <=  std_logic_vector(unsigned(var) ror 22);
					elsif(Cs = "10110") then
						v1 <=  std_logic_vector(unsigned(var) ror 23);
					elsif(Cs = "10111") then
						v1 <=  std_logic_vector(unsigned(var) ror 24);
					elsif(Cs = "11000") then
						v1 <=  std_logic_vector(unsigned(var) ror 25);
					elsif(Cs = "11001") then
						v1 <=  std_logic_vector(unsigned(var) ror 25);
					elsif(Cs = "11010") then
						v1 <=  std_logic_vector(unsigned(var) ror 26);
					elsif(Cs = "11011") then
						v1 <=  std_logic_vector(unsigned(var) ror 27);
					elsif(Cs = "11100") then
						v1 <=  std_logic_vector(unsigned(var) ror 28);
					elsif(Cs = "11101") then
						v1 <=  std_logic_vector(unsigned(var) ror 29);
					elsif(Cs = "11110") then
						v1 <=  std_logic_vector(unsigned(var) ror 30);
					elsif(Cs = "11111") then
						v1 <=  std_logic_vector(unsigned(var) ror 31);
					end if;
			end if;		
	end process;
	Sout <= v1;
end beh;
